library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity ROM_16_8 IS
	port(address : in std_logic_vector(3 downto 0);
			dataOut : out std_logic_vector(7 downto 0));
end ROM_16_8;

architecture Behav of ROM_16_8 is
	
	subtype Dataword is std_logic_vector(7 downto 0);
	type TROM is array (0 to 15) of Dataword;
	
constant ROMcontent : TROM := (X"01",X"02",X"04",X"08",
										 X"03",X"06",X"0C",X"18",
										 X"07",X"0E",X"1C",X"38",
										 X"0F",X"1E",X"3C",X"78");

begin
	
	dataOut <= ROMcontent(to_integer(unsigned(address)));
	
end Behav;