-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 17.1.0 Build 590 10/25/2017 SJ Lite Edition
-- Created on Thu May 16 09:44:50 2019

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY DrinksFSM IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        m20 : IN STD_LOGIC := '0';
        m50 : IN STD_LOGIC := '0';
        drink : OUT STD_LOGIC
    );
END DrinksFSM;

ARCHITECTURE BEHAVIOR OF DrinksFSM IS
    TYPE type_fstate IS (ST0,ST1,ST2,ST3,ST4,ST5);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,m20,m50)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= ST0;
            drink <= '0';
        ELSE
            drink <= '0';
            CASE fstate IS
                WHEN ST0 =>
                    IF (((m20 = '0') AND (m50 = '0'))) THEN
                        reg_fstate <= ST0;
                    ELSIF (((m20 = '1') AND (m50 = '0'))) THEN
                        reg_fstate <= ST1;
                    ELSIF (((m20 = '0') AND (m50 = '1'))) THEN
                        reg_fstate <= ST2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ST0;
                    END IF;

                    drink <= '0';
                WHEN ST1 =>
                    IF (((m20 = '0') AND (m50 = '0'))) THEN
                        reg_fstate <= ST1;
                    ELSIF (((m20 = '1') AND (m50 = '0'))) THEN
                        reg_fstate <= ST2;
                    ELSIF (((m20 = '0') AND (m50 = '1'))) THEN
                        reg_fstate <= ST3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ST1;
                    END IF;

                    drink <= '0';
                WHEN ST2 =>
                    IF (((m20 = '0') AND (m50 = '0'))) THEN
                        reg_fstate <= ST2;
                    ELSIF (((m20 = '1') AND (m50 = '0'))) THEN
                        reg_fstate <= ST3;
                    ELSIF (((m20 = '0') AND (m50 = '1'))) THEN
                        reg_fstate <= ST4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ST2;
                    END IF;

                    drink <= '0';
                WHEN ST3 =>
                    IF (((m20 = '0') AND (m50 = '0'))) THEN
                        reg_fstate <= ST3;
                    ELSIF (((m20 = '1') AND (m50 = '0'))) THEN
                        reg_fstate <= ST4;
                    ELSIF (((m20 = '0') AND (m50 = '1'))) THEN
                        reg_fstate <= ST5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ST3;
                    END IF;

                    drink <= '0';
                WHEN ST4 =>
                    IF (((m20 = '0') AND (m50 = '0'))) THEN
                        reg_fstate <= ST4;
                    ELSIF (((m20 = '1') OR (m50 = '1'))) THEN
                        reg_fstate <= ST5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ST4;
                    END IF;

                    drink <= '0';
                WHEN ST5 =>
                    IF (((m20 = '0') AND (m50 = '0'))) THEN
                        reg_fstate <= ST0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ST5;
                    END IF;

                    drink <= '1';
                WHEN OTHERS => 
                    drink <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
